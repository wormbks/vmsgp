module vmsgp
