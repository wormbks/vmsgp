module msgp
