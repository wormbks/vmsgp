module msgp

//{	"string": "foo bar" }
const foo_bar_as_map = [u8(0x81), 0xA6, 0x73, 0x74, 0x72, 0x69, 0x6E, 0x67, 0xA7, 0x66, 0x6F, 0x6F,
	0x20, 0x62, 0x61, 0x72] // this one is map

const foo_bar_as_tuple = [u8(0xA6), 0x73, 0x74, 0x72, 0x69, 0x6E, 0x67, 0xA7, 0x66, 0x6F, 0x6F,
	0x20, 0x62, 0x61, 0x72]

fn test_read_string_len() {
	mut br := BufReader{
		buf: foo_bar_as_tuple
		len: foo_bar_as_tuple.len
	}
	mut s := Decoder{
		br: br
	}
	l := s.string_length() or { 0 }
	assert l == 6
}

fn test_read_string() {
	mut br := BufReader{
		buf: foo_bar_as_tuple
		len: foo_bar_as_tuple.len
	}
	mut s := Decoder{
		br: br
	}
	l := s.read_string() or { '' }
	assert l.len == 6
}

fn write_fix_sring() {
	str := '1234567890' //[u8(0xAA), 0x30, 0x31, 0x32, 0x33, 0x34, 0x35, 0x36, 0x37, 0x38, 0x39]
	mut bw := make_buf_writer(str.len + 2)
	mut w := Encoder{
		bw: bw
	}
	w.write_sring(str) or { -1 }
	assert bw.buf[0] == 0xAA
	assert bw.buf[3] == 0x32
}

fn write_short_sring() {
	str := '0123456789012345678901234567890123456789'
	// 0xD9, 0x28, 0x30, 0x31, 0x32, 0x33, 0x34, 0x35, 0x36, 0x37, 0x38, 0x39, 0x30, 0x31, 0x32, 0x33, 0x34, 0x35, 0x36, 0x37, 0x38, 0x39, 0x30, 0x31, 0x32, 0x33, 0x34, 0x35, 0x36, 0x37, 0x38, 0x39, 0x30, 0x31, 0x32, 0x33, 0x34, 0x35, 0x36, 0x37, 0x38, 0x39
	mut bw := make_buf_writer(str.len + 2)
	mut w := Encoder{
		bw: bw
	}
	w.write_sring(str) or { -1 }
	assert bw.buf[0] == 0xD9
	assert bw.buf[1] == 0x28
	assert bw.buf[2] == 0x30
	assert bw.buf[3] == 0x30
}
